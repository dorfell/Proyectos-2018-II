library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package phrases is

type palabra_1 is array ( 0 to 80) of std_logic_vector (7 downto 0);
type palabra_2 is array ( 0 to 36) of std_logic_vector (7 downto 0);
type palabra_3 is array ( 0 to 60) of std_logic_vector (7 downto 0);
type palabra_4 is array ( 0 to 113) of std_logic_vector (7 downto 0);
type palabra_5 is array ( 0 to 169) of std_logic_vector (7 downto 0);
type palabra_6 is array ( 0 to 28) of std_logic_vector (7 downto 0);
type palabra_7 is array ( 0 to 210) of std_logic_vector (7 downto 0);

constant w_id : palabra_1;
constant w_sent : palabra_2;
constant w_code : palabra_3;
constant w_question : palabra_4;
constant w_finish : palabra_5;
constant w_error : palabra_6;
constant w_check : palabra_7;

end phrases;

package body phrases is

constant w_id : palabra_1 := ( 
"01111111","01000001","01000001","01000001","00111110","00000000", --D
"00101111","00000000", --i
"00011000","00100101","00100101","00100101","00011110","00000000", --g
"00101111","00000000", --i
"00010000","01111111","00010000","00000000", --t
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00000000","00000000","00000000", --espacio
"00001110","00010001","00010001","00010001","01111111","00000000", --d
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00001110","00010001","00010001","00010001","00010001","00000000", --c
"00011110","00000001","00000001","00000001","00011110","00000000", --u
"00011111","00010000","00001100","00010000","00011111","00000000", --m
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00011111","00001000","00010000","00010000","00011111","00000000", --n
"00010000","01111111","00010000","00000000", --t
"00001110","00010001","00010001","00010001","00001110","00000000" --o
); --81

constant w_sent : palabra_2 := (
"01111111","01001001","01001001","01001001","01000001","00000000", --E
"00011111","00001000","00010000","00010000","00011111","00000000", --n
"00011100","00000010","00000001","00000010","00011100","00000000", --v
"00101111","00000000", --i
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00001110","00010001","00010001","00010001","01111111","00000000", --d
"00001110","00010001","00010001","00010001","00001110" --o
); --37

constant w_code : palabra_3 := ( 
"01111111","01000001","01000001","01000001","00111110","00000000", --D
"00101111","00000000", --i
"00011000","00100101","00100101","00100101","00011110","00000000", --g
"00101111","00000000", --i
"00010000","01111111","00010000","00000000", --t
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00000000","00000000","00000000", --espacio
"00001110","00010001","00010001","00010001","00010001","00000000", --c
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00001110","00010001","00010001","00010001","01111111","00000000", --d
"00101111","00000000", --i
"00011000","00100101","00100101","00100101","00011110","00000000", --g
"00001110","00010001","00010001","00010001","00001110","00000000" --o
); --61

constant w_question : palabra_4 := ( 
"00000110","00001001","01010001","00000001","00000010","00000000", --�
"00110010","01001001","01001001","01001001","00100110","00000000", --S
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00011000","00100101","00100101","00100101","00011110","00000000", --g
"00011110","00000001","00000001","00000001","00011110","00000000", --u
"00101111","00000000", --i
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00000000","00000000","00000000", --espacio
"00001110","00010001","00010001","00010001","00010001","00000000", --c
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00011111","00001000","00010000","00010000","00011111","00000000", --n
"00000000","00000000","00000000", --espacio
"00011111","00100100","00100100","00100100","00011000","00000000", --p
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00001001","00010101","00010101","00010101","00010010","00000000", --s
"00010000","01111111","00010000","00000000", --t
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00011111","00010000","00001100","00010000","00011111","00000000", --m
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00100000","01000000","01001101","01010000","00100000","00000000" --?
); --114

constant w_finish : palabra_5 := ( 
"01111111","01001000","01001000","01001000","00110000","00000000", --P
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00001001","00010101","00010101","00010101","00010010","00000000", --s
"00010000","01111111","00010000","00000000", --t
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00011111","00010000","00001100","00010000","00011111","00000000", --m
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00000000","00000000","00000000", --espacio
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"01111111","00000000", --l
"00101111","00000000", --i
"00010001","00010011","00010101","00011001","00010001","00000000", --z
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00001110","00010001","00010001","00010001","01111111","00000000", --d
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00001101","00001110","00000000", --,
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00001001","00010101","00010101","00010101","00010010","00000000", --s
"00011111","00100100","00100100","00100100","00011000","00000000", --p
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00000000","00000000","00000000", --espacio
"01111111","00000000", --l
"01111111","00000000", --l
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00011111","00010000","00001100","00010000","00011111","00000000", --m
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00001110","00010001","00010001","00010001","01111111","00000000", --d
"00001110","00010001","00010001","00010001","00001110" --o
); --170

constant w_error : palabra_6 := ( 
"01111111","01001001","01001001","01001001","01000001","00000000", --E
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010001","00010001","00010001","00001110", --o
"00010000","00001111","00010000","00010000","00010000","00000000" --r
); --29

constant w_check : palabra_7 := ( 
"01111111","01001001","01001001","01001001","01000001","00000000", --E
"00011111","00001000","00010000","00010000","00011111","00000000", --n
"00010000","01111111","00010000","00000000", --t
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00000000","00000000","00000000", --espacio
"00011111","00100100","00100100","00100100","00011000","00000000", --p
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00000000","00000000","00000000", --espacio
"00001110","00010001","00010001","00010001","00010001","00000000", --c
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00011111","00001000","00010000","00010000","00011111","00000000", --n
"00001000","00111111","01001000","00100000","00000000", --f
"00101111","00000000", --i
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00011111","00010000","00001100","00010000","00011111","00000000", --m
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00000000","00000000","00000000", --espacio
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00000000","00000000","00000000", --espacio
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00001001","00010101","00010101","00010101","00010010","00000000", --s
"00001110","00010001","00010001","00010001","00010001","00000000", --c
"00000000","00000000","00000000", --espacio
"00011111","00100100","00100100","00100100","00011000","00000000", --p
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010001","00010001","00011111","00000001","00000000", --a
"00000000","00000000","00000000", --espacio
"00001110","00010001","00010001","00010001","00010001","00000000", --c
"00001110","00010001","00010001","00010001","00001110","00000000", --o
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00010000","00001111","00010000","00010000","00010000","00000000", --r
"00001110","00010101","00010101","00010101","00001000","00000000", --e
"00011000","00100101","00100101","00100101","00011110","00000000", --g
"00101111","00000000", --i
"00010000","00001111","00010000","00010000","00010000","00000000" --r
); --211

end package body phrases;

--A => "00111111","01001000","01001000","01001000","00111111"
--B => "01111111","01001001","01001001","01001001","00110110"
--C => "00111110","01000001","01000001","01000001","00100010"
--D => "01111111","01000001","01000001","01000001","00111110"
--E => "01111111","01001001","01001001","01001001","01000001"
--F => "01111111","01001000","01001000","01001000","01000000"
--G => "01111110","01000001","01001001","01001001","00101110"
--H => "01111111","00001000","00001000","00001000","01111111"
--I => "01000001","01111111","01000001"
--J => "00000010","00000001","00000001","00000001","01111110"
--K => "01111111","00001000","00010100","00100010","01000001"
--L => "01111111","00000001","00000001","00000001","00000001"
--M => "01111111","00100000","00010000","00100000","01111111"
--N => "01111111","00010000","00001000","00000100","01111111"
--� => "01111111","10010000","10001000","10000100","01111111"
--O => "00111110","01000001","01000001","01000001","00111110"
--P => "01111111","01001000","01001000","01001000","00110000"
--Q => "00111110","01000001","01000101","01000011","00111111"
--R => "01111111","01001000","01001100","01001010","00110001"
--S => "00110010","01001001","01001001","01001001","00100110"
--T => "01000000","01000000","01111111","01000000","01000000"
--U => "01111110","00000001","00000001","00000001","01111110"
--V => "01111100","00000010","00000001","00000010","01111100"
--W => "01111111","00000010","00000100","00000010","01111110"
--X => "01100011","00010100","00001000","00010100","01100011"
--Y => "01110000","00001000","00000111","00001000","01110000"
--Z => "01000011","01000101","01001001","01010001","01100001"

--a => "00001110","00010001","00010001","00011111","00000001"
--b => "01111111","00010001","00010001","00010001","00001110"
--c => "00001110","00010001","00010001","00010001","00001010"
--d => "00001110","00010001","00010001","00010001","01111111"
--e => "00001110","00010101","00010101","00010101","00001000"
--f => "00001000","00111111","01001000","00100000"
--g => "00011000","00100101","00100101","00100101","00011110"
--h => "01111111","00010000","00010000","00010000","00001111"
--i => "01011111"
--j => "00000010","00000001","00000001","01011110"
--k => "01111111","00000100","00000100","00001010","00010001"
--l => "01111111"
--m => "00011111","00010000","00001100","00010000","00011111"
--n => "00011111","00001000","00010000","00010000","00011111"
--� => "00011111","01001000","01010000","01010000","00011111"
--o => "00001110","00010001","00010001","00010001","00001110"
--p => "00011111","00100100","00100100","00100100","00011000"
--q => "00011000","00100100","00100100","00100100","00011111"
--r => "00010000","00001111","00010000","00010000","00010000",
--s => "00001001","00010101","00010101","00010101","00010010"
--t => "00010000","01111111","00100000"
--u => "00011110","00000001","00000001","00000001","00011110"
--v => "00011100","00000010","00000001","00000010","00011100"
--w => "00011110","00000001","00000110","00000001","00011110"
--x => "00010001","00001010","00000100","00001010","00010001"
--y => "00010000","00001000","00000111","00001000","00010000"
--z => "00010001","00010011","00010101","00011001","00010001"

--0 => "00111110","01000101","01001001","01010001","00111110"
--1 => "00100001","01111111","00000001" 
--2 => "00100001","01000011","01000101","01001001","00110001"
--3 => "00100010","01000001","01001001","01001001","00110110"
--4 => "00000100","00001100","00010100","00100100","01111111"
--5 => "01111001","01001001","01001001","01001001","01000110"
--6 => "00111110","01001001","01001001","01001001","00100110"
--7 => "01000000","01000000","01000111","01001000","01110000"
--8 => "00110110","01001001","01001001","01001001","00110110"
--9 => "00110010","01001001","01001001","01001001","00111110"

--� => "00100000","01010000","01001101","01000000","00100000"
--? => "00100000","01000000","01001101","01010000","00100000"
--, => "00001101","00001110"
