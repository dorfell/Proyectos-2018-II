-- contador mod m para el módulo UART
-- Baudrate 9600;
-- Sampling ticks 32;
-- reloj 50MHz;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mcounter is
	generic (
		N: integer := 8;   -- 8 bits para llega a 256
		M: integer := 163 -- 163 modulo para UART
	);
	port (
		clk, reset: in	std_logic;
		max_tick: out std_logic;
		q: out	std_logic_vector (N-1 downto 0)
	);
end mcounter;

architecture Behavioral of mcounter is
	signal r_reg, r_next: unsigned (N-1 downto 0);

begin
	-- registro
	process (clk,reset)
	begin
		if (reset = '1') then
			r_reg <= (others =>'0');
		elsif (clk'event and clk='1') then
			r_reg <= r_next;
		end if;
	end process;
	
	-- lógica
	r_next <= (others => '0') when r_reg = (M-1) else r_reg + 1;
	
	-- salida
	q <= std_logic_vector(r_reg);
	max_tick <= '1' when r_reg = (M-1) else '0';
end Behavioral;